`ifndef PULPINO_SPI_MASTER_SUBSYSTEM_VIRTUAL_SEQ_PKG_INCLUDED_
`define PULPINO_SPI_MASTER_SUBSYSTEM_VIRTUAL_SEQ_PKG_INCLUDED_

//--------------------------------------------------------------------------------------------
// Package : pulpino_spi_master_subsystem_virtual_seq_pkg
// Includes all the master seq files declared
//--------------------------------------------------------------------------------------------
package pulpino_spi_master_subsystem_virtual_seq_pkg;

  //-------------------------------------------------------
  // Importing UVM Pkg
  //-------------------------------------------------------
  `include "uvm_macros.svh"
  import uvm_pkg::*;

  import axi4_master_pkg::*;
  import spi_slave_pkg::*;
  import axi4_master_seq_pkg::*;
  import spi_slave_seq_pkg::*;
  import env_pkg::*;
  import axi4_reg_seq_pkg::*;

  //-------------------------------------------------------
  // Including required package files
  //-------------------------------------------------------
  `include "virtual_base_seq.sv"
  `include "virtual_basic_write_read_reg_seq.sv"
  `include "virtual_basic_write_seq.sv"
  `include "virtual_basic_read_seq.sv"
  
  // Register virtual sequences
  `include "virtual_reg_seq.sv"
  `include "virtual_std_mode_write_0_cmd_0_addr_32_data_length_reg_seq.sv"
  `include "virtual_std_mode_write_0_cmd_0_addr_16_data_length_reg_seq.sv"
  `include "virtual_std_mode_write_0_cmd_16_addr_16_data_length_reg_seq.sv"
  `include "virtual_std_mode_write_16_cmd_16_addr_16_data_length_reg_seq.sv"
  `include "virtual_std_mode_write_0_cmd_32_addr_32_data_length_reg_seq.sv"
  `include "virtual_std_mode_write_32_cmd_32_addr_32_data_length_reg_seq.sv"

  `include "virtual_std_mode_write_16_cmd_16_addr_32_data_length_reg_seq.sv"
  `include "virtual_std_mode_write_8_cmd_32_addr_32_data_length_reg_seq.sv"
  `include "virtual_std_mode_write_8_cmd_8_addr_32_data_length_reg_seq.sv"
  `include "virtual_std_mode_write_8_cmd_16_addr_32_data_length_reg_seq.sv"
  `include "virtual_std_mode_write_even_clkdiv_reg_seq.sv"

  `include "virtual_spi_modes_clkdiv_dummy_cycles_cross_reg_seq.sv"
  `include "virtual_spi_modes_transfer_length_interupts_cross_reg_seq.sv"

  //`include "virtual_rand_reg_seq.sv"


endpackage : pulpino_spi_master_subsystem_virtual_seq_pkg

`endif
