`ifndef PULPINO_SPI_MASTER_SUBSYSTEM_VIRTUAL_BASIC_WRITE_READ_REG_SEQ_INCLUDED_
`define PULPINO_SPI_MASTER_SUBSYSTEM_VIRTUAL_BASIC_WRITE_READ_REG_SEQ_INCLUDED_

//--------------------------------------------------------------------------------------------
// Class: pulpino_spi_master_subsystem_virtual_basic_write_read_reg_seq
// <Descrsubsystemtion_here>
//--------------------------------------------------------------------------------------------
class pulpino_spi_master_subsystem_virtual_basic_write_read_reg_seq extends pulpino_spi_master_subsystem_virtual_base_seq;
  `uvm_object_utils(pulpino_spi_master_subsystem_virtual_basic_write_read_reg_seq)

  axi4_master_basic_write_read_reg_seq axi4_master_basic_write_read_reg_seq_h;
  spi_fd_basic_slave_seq spi_fd_basic_slave_seq_h;

  //Variable : write_read_key
  //Used to provide access to perform write and read operation
  semaphore write_read_key;

  

  //-------------------------------------------------------
  // Externally defined Tasks and Functions
  //-------------------------------------------------------
  extern function new(string name = "pulpino_spi_master_subsystem_virtual_basic_write_read_reg_seq");
  extern task body();
endclass : pulpino_spi_master_subsystem_virtual_basic_write_read_reg_seq

//--------------------------------------------------------------------------------------------
// Construct: new
//
// Parameters:
//  name - pulpino_spi_master_subsystem_virtual_basic_write_read_reg_seq
//--------------------------------------------------------------------------------------------
function pulpino_spi_master_subsystem_virtual_basic_write_read_reg_seq::new(string name = "pulpino_spi_master_subsystem_virtual_basic_write_read_reg_seq");
  super.new(name);
  write_read_key = new(1);
endfunction : new

//--------------------------------------------------------------------------------------------
// Task - body
// Creates a master reqister sequence and slave normal sequence
//--------------------------------------------------------------------------------------------
task pulpino_spi_master_subsystem_virtual_basic_write_read_reg_seq::body();
  super.body();

  fork
    forever begin : SLAVE_SEQ
      `uvm_info("slave_vseq",$sformatf("started slave vseq"),UVM_HIGH)
      write_read_key.get(1);
      spi_fd_basic_slave_seq_h = spi_fd_basic_slave_seq::type_id::create("spi_fd_basic_slave_seq_h");
      spi_fd_basic_slave_seq_h.start(p_sequencer.spi_slave_seqr_h);
      write_read_key.put(1);
      `uvm_info("slave_vseq",$sformatf("ended slave vseq"),UVM_HIGH)
    end
  join_none

  repeat(1) begin
   `uvm_info("master_vseq",$sformatf("started master vseq"),UVM_HIGH)
   write_read_key.get(1);
   axi4_master_basic_write_read_reg_seq_h = axi4_master_basic_write_read_reg_seq::type_id::create("axi4_master_basic_write_read_reg_seq_h");
   axi4_master_basic_write_read_reg_seq_h.model = p_sequencer.env_config_h.spi_master_reg_block;
   axi4_master_basic_write_read_reg_seq_h.start(p_sequencer.axi4_master_write_seqr_h);
   //axi4_master_basic_write_read_reg_seq_h.start(p_sequencer.axi4_master_read_seqr_h);
   write_read_key.put(1);
   `uvm_info("master_vseq",$sformatf("ended master vseq"),UVM_HIGH)
 end
 endtask : body


`endif
